** Profile: "SCHEMATIC1-siim1"  [ C:\Users\asus\Desktop\New folder\p1-pspicefiles\schematic1\siim1.sim ] 

** Creating circuit file "siim1.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "C:/Cadence/SPB_17.2/tools/capture/library/pspice/BC846B.lib" 
* From [PSPICE NETLIST] section of C:\Users\asus\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
